`include "controller.v"
`timescale 1ns / 1ps

module controller_tb;

// Declaración de señales del controlador
reg clk, reset;
// Otras señales del controlador...

// Instancia del módulo controlador
controller_instance controller_inst (
    .clk(clk),
    .reset(reset),
    // Otras señales del controlador...
);

// Inicialización de señales
initial begin
    $dumpfile("controller/sim.vcd");
    $dumpvars(0, controller_tb);

    clk = 0;
    reset = 1;
    // Inicialización de otras señales...

    // Generación de estímulos para el controlador...
end

// Generación de reloj
always #5 clk = ~clk;

endmodule