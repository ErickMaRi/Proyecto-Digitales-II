module peripheral(
    input clk,
    input reset)
;

endmodule